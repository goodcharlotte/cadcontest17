module WHY ( g7 , g29 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 , g119 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 , t_0 , g30 , g41 , g51 , g62 , g124 , g217 , g_g217 );
input g7 , g29 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 , g119 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 , t_0 , g30 , g41 , g51 , g62 , g124 ;
output g217 , g_g217 ;
wire n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , g_g217 , g_n80 , g_n81 , g_n82 , g_n83 , g_n84 , g_n85 , g_n86 , g_n87 , g_n88 , g_n89 , g_n90 , g_n91 , g_n92 , g_n93 , g_n94 , g_n95 , g_n96 , g_n97 , g_n98 , g_n99 , g_n100 , g_n101 , g_n102 , g_n103 , g_n104 , g_n105 , g_n106 , g_n107 , g_n108 , g_n109 , g_n110 , g_n111 , g_n112 , g_n113 , g_n114 , g_n115 , g_n116 , g_n117 , g_n118 , g_n119 , g_n120 , g_n121 , g_n122 , g_n123 , g_n124 , g_n125 , g_n126 , g_n127 , g_n128 , g_n129 , g_n130 , g_n131 , g_n132 , g_n133 , g_n134 , g_n135 , g_n136 , g_n137 , g_n138 , g_n139 , g_n140 , g_n141 , g_n142 , g_n143 , g_n144 , g_n145 , g_n146 , g_n147 , g_n148 , g_n149 , g_n150 , g_n151 , g_n152 , g_n153 , g_n154 , g_n155 , g_n156 , g_n157 , g_n158 , g_n159 , g_n160 , g_n161 , g_n162 , g_n163 , g_n164 , g_n165 , g_n166 , g_n167 , g_n168 , g_n169 , g_n170 , g_n171 , g_n172 , g_n173 , g_n174 , g_n175 , g_n176 , g_n177 , g_n178 , g_n179 , g_n180 , g_n181 , g_n182 , g_n183 , g_n184 , g_n185 , g_n186 , g_n187 , g_n188 , g_n189 , g_n190 , g_n191 , g_n192 , g_n193 , g_n194 , g_n195 , g_n196 , g_n197 , g_n198 , g_n199 , g_n200 , g_n201 , g_n202 , g_n203 , g_n204 , g_n205 , g_n206 , g_n207 , g_n208 , g_n209 , g_n210 , g_n211 , g_n212 , g_n213 , g_n214 , g_n215 , g_n216 , g_n217 , g_n218 , g_n219 , g_n220 , g_n221 , g_n222 , g_n223 , g_n224 , g_n225 , g_n226 , g_n227 , g_n228 , g_n229 , g_n230 , g_n231 , g_n232 , g_n233 , g_n234 , g_n235 , g_n236 , g_n237 , g_n238 , g_n239 , g_n240 , g_n241 , g_n242 , g_n243 , g_n244 , g_n245 , g_n246 , g_n247 , g_n248 , g_n249 , g_n250 , g_n251 , g_n252 , g_n253 , g_n254 , g_n255 , g_n256 , g_n257 , g_n258 , g_n259 , g_n260 , g_n261 , g_n262 , g_n263 , g_n264 , g_n265 , g_n266 , g_n267 , g_n268 , g_n269 , g_n270 , g_n271 , g_n272 , g_n273 , g_n274 , g_n275 , g_n276 , g_n277 , g_n278 , g_n279 , g_n280 , g_n281 , g_n282 , g_n283 , g_n284 , g_n285 , g_n286 , g_n287 , g_n288 , g_n289 , g_n290 , g_n291 , g_n292 , g_n293 , g_n294 ;
nor ( n80 , g116 , g46 );
or ( n81 , n80 , n79 );
or ( n82 , n81 , n78 );
nor ( n83 , n77 , g36 );
nor ( n84 , g116 , g68 );
or ( n85 , n84 , g119 );
or ( n86 , n85 , n83 );
and ( n87 , n86 , n82 );
or ( n88 , n87 , n76 );
nor ( n89 , n79 , g58 );
nor ( n90 , g119 , g37 );
or ( n91 , n90 , n77 );
or ( n92 , n91 , n89 );
nor ( n93 , n79 , g47 );
nor ( n94 , g119 , g69 );
or ( n95 , n94 , g116 );
or ( n96 , n95 , n93 );
and ( n97 , n96 , n92 );
not ( n98 , g144 );
and ( n99 , g145 , n98 );
and ( n100 , n99 , g99 );
not ( n101 , g145 );
and ( n102 , n101 , g144 );
and ( n103 , n102 , g79 );
nor ( n104 , n103 , n100 );
and ( n105 , g145 , g144 );
and ( n106 , n105 , g89 );
and ( n107 , n101 , n98 );
and ( n108 , n107 , g109 );
nor ( n109 , n108 , n106 );
and ( n110 , n109 , n104 );
nor ( n111 , n110 , g126 );
and ( n112 , n102 , g78 );
not ( n113 , n112 );
and ( n114 , n113 , g29 );
and ( n115 , n99 , g98 );
not ( n116 , n115 );
and ( n117 , n107 , g108 );
and ( n118 , n105 , g88 );
nor ( n119 , n118 , n117 );
and ( n120 , n119 , n116 );
and ( n121 , n120 , n114 );
and ( n122 , n121 , n111 );
not ( n123 , n122 );
nand ( n124 , n123 , g128 );
nand ( n125 , n122 , g139 );
and ( n126 , n125 , n124 );
or ( n127 , n126 , n97 );
and ( n128 , n126 , n97 );
nor ( n129 , n77 , g59 );
nor ( n130 , g116 , g48 );
or ( n131 , n130 , n79 );
or ( n132 , n131 , n129 );
nor ( n133 , n77 , g38 );
nor ( n134 , g116 , g70 );
or ( n135 , n134 , g119 );
or ( n136 , n135 , n133 );
and ( n137 , n136 , n132 );
nand ( n138 , n123 , g127 );
nand ( n139 , n122 , g138 );
and ( n140 , n139 , n138 );
or ( n141 , n140 , n137 );
and ( n142 , n140 , n137 );
nor ( n143 , n77 , g60 );
nor ( n144 , g116 , g49 );
or ( n145 , n144 , n79 );
or ( n146 , n145 , n143 );
nor ( n147 , n77 , g39 );
nor ( n148 , g116 , g71 );
or ( n149 , n148 , g119 );
or ( n150 , n149 , n147 );
and ( n151 , n150 , n146 );
or ( n152 , n151 , t_0 );
and ( n153 , n151 , t_0 );
nand ( n154 , n123 , g125 );
not ( n155 , g137 );
or ( n156 , n123 , n155 );
and ( n157 , n156 , n154 );
or ( n158 , n157 , n153 );
and ( n159 , n158 , n152 );
or ( n160 , n159 , n142 );
and ( n161 , n160 , n141 );
or ( n162 , n161 , n128 );
and ( n163 , n162 , n127 );
or ( n164 , n163 , n88 );
nand ( n165 , n123 , g129 );
nand ( n166 , n122 , g140 );
and ( n167 , n166 , g7 );
and ( n168 , n167 , n165 );
and ( n169 , n168 , n164 );
nor ( n170 , n77 , g56 );
nor ( n171 , g116 , g45 );
or ( n172 , n171 , n79 );
or ( n173 , n172 , n170 );
nor ( n174 , n77 , g35 );
nor ( n175 , g116 , g67 );
or ( n176 , n175 , g119 );
or ( n177 , n176 , n174 );
and ( n178 , n177 , n173 );
or ( n179 , n178 , n76 );
nand ( n180 , n123 , g130 );
nand ( n181 , n122 , g141 );
and ( n182 , n181 , g7 );
and ( n183 , n182 , n180 );
and ( n184 , n183 , n179 );
and ( n185 , n163 , n88 );
or ( n186 , n185 , n184 );
or ( n187 , n186 , n169 );
or ( n188 , n183 , n179 );
and ( n189 , n123 , g7 );
not ( n190 , n189 );
and ( n191 , g119 , g55 );
not ( n192 , n191 );
and ( n193 , n79 , g34 );
nor ( n194 , n193 , n77 );
and ( n195 , n194 , n192 );
nor ( n196 , g116 , g66 );
and ( n197 , n196 , n79 );
nor ( n198 , n197 , n195 );
xor ( n199 , n198 , g131 );
or ( n200 , n199 , n190 );
not ( n201 , g132 );
nor ( n202 , n77 , g54 );
not ( n203 , n202 );
nor ( n204 , g116 , g44 );
nor ( n205 , n204 , n79 );
and ( n206 , n205 , n203 );
nor ( n207 , n77 , g33 );
not ( n208 , n207 );
nor ( n209 , g116 , g65 );
nor ( n210 , n209 , g119 );
and ( n211 , n210 , n208 );
nor ( n212 , n211 , n206 );
or ( n213 , n212 , n201 );
or ( n214 , n213 , n190 );
and ( n215 , n212 , n201 );
and ( n216 , n215 , n189 );
not ( n217 , n216 );
and ( n218 , n217 , n214 );
and ( n219 , n218 , n200 );
and ( n220 , n219 , n188 );
and ( n221 , n220 , n187 );
nor ( n222 , n198 , g131 );
and ( n223 , n222 , n189 );
and ( n224 , n223 , n214 );
or ( n225 , n224 , n216 );
or ( n226 , n225 , n221 );
not ( n227 , n111 );
and ( n228 , n121 , n227 );
not ( n229 , n228 );
and ( n230 , n102 , g81 );
and ( n231 , n105 , g91 );
nor ( n232 , n231 , n230 );
and ( n233 , n107 , g111 );
and ( n234 , n99 , g101 );
nor ( n235 , n234 , n233 );
and ( n236 , n235 , n232 );
nor ( n237 , n236 , n229 );
not ( n238 , n237 );
or ( n239 , n238 , n155 );
and ( n240 , n228 , n155 );
and ( n241 , n240 , n238 );
not ( n242 , n241 );
and ( n243 , n242 , n239 );
not ( n244 , g134 );
and ( n245 , n99 , g94 );
and ( n246 , n105 , g84 );
nor ( n247 , n246 , n245 );
and ( n248 , n102 , g74 );
and ( n249 , n107 , g104 );
nor ( n250 , n249 , n248 );
and ( n251 , n250 , n247 );
or ( n252 , n251 , n244 );
nor ( n253 , n252 , n229 );
and ( n254 , n251 , n244 );
and ( n255 , n254 , n228 );
nor ( n256 , n255 , n253 );
and ( n257 , n256 , n243 );
and ( n258 , n99 , g102 );
and ( n259 , n105 , g92 );
nor ( n260 , n259 , n258 );
and ( n261 , n102 , g82 );
and ( n262 , n107 , g112 );
nor ( n263 , n262 , n261 );
and ( n264 , n263 , n260 );
nor ( n265 , n264 , n229 );
and ( n266 , n265 , g135 );
not ( n267 , n265 );
nor ( n268 , n229 , g135 );
and ( n269 , n268 , n267 );
nor ( n270 , n269 , n266 );
not ( n271 , g133 );
nor ( n272 , n77 , g53 );
not ( n273 , n272 );
nor ( n274 , g116 , g43 );
nor ( n275 , n274 , n79 );
and ( n276 , n275 , n273 );
nor ( n277 , n77 , g32 );
not ( n278 , n277 );
nor ( n279 , g116 , g64 );
nor ( n280 , n279 , g119 );
and ( n281 , n280 , n278 );
nor ( n282 , n281 , n276 );
and ( n283 , n282 , n271 );
and ( n284 , n283 , n228 );
or ( n285 , n282 , n271 );
nor ( n286 , n285 , n229 );
nor ( n287 , n286 , n284 );
and ( n288 , n287 , n270 );
and ( n289 , n288 , n257 );
and ( n290 , n289 , n226 );
and ( n291 , n255 , n243 );
and ( n292 , n291 , n270 );
and ( n293 , n284 , n270 );
and ( n294 , n293 , n257 );
and ( n295 , n269 , n239 );
or ( n296 , n295 , n241 );
or ( n297 , n296 , n294 );
or ( n298 , n297 , n292 );
or ( g_g217 , g_n294 , g_n282 );
and ( g_n80 , g145 , g88 );
not ( g_n81 , g_n80 );
not ( g_n82 , g144 );
not ( g_n83 , g145 );
and ( g_n84 , g_n83 , g78 );
nor ( g_n85 , g_n84 , g_n82 );
and ( g_n86 , g_n85 , g_n81 );
and ( g_n87 , g145 , g98 );
not ( g_n88 , g_n87 );
and ( g_n89 , g_n83 , g108 );
nor ( g_n90 , g_n89 , g144 );
and ( g_n91 , g_n90 , g_n88 );
nor ( g_n92 , g_n91 , g_n86 );
not ( g_n93 , g_n92 );
and ( g_n94 , g_n93 , g29 );
nor ( g_n95 , g_n83 , g89 );
not ( g_n96 , g_n95 );
nor ( g_n97 , g145 , g79 );
nor ( g_n98 , g_n97 , g_n82 );
and ( g_n99 , g_n98 , g_n96 );
nor ( g_n100 , g_n83 , g99 );
not ( g_n101 , g_n100 );
nor ( g_n102 , g145 , g109 );
nor ( g_n103 , g_n102 , g144 );
and ( g_n104 , g_n103 , g_n101 );
nor ( g_n105 , g_n104 , g_n99 );
nor ( g_n106 , g_n105 , g126 );
not ( g_n107 , g_n106 );
and ( g_n108 , g_n107 , g_n94 );
not ( g_n109 , g_n108 );
not ( g_n110 , g135 );
nand ( g_n111 , g144 , g92 );
nand ( g_n112 , g_n82 , g102 );
and ( g_n113 , g_n112 , g145 );
and ( g_n114 , g_n113 , g_n111 );
nand ( g_n115 , g144 , g82 );
nand ( g_n116 , g_n82 , g112 );
and ( g_n117 , g_n116 , g_n83 );
and ( g_n118 , g_n117 , g_n115 );
or ( g_n119 , g_n118 , g_n114 );
or ( g_n120 , g_n119 , g_n110 );
not ( g_n121 , g133 );
not ( g_n122 , g116 );
not ( g_n123 , g119 );
and ( g_n124 , g_n123 , g_n122 );
nand ( g_n125 , g_n124 , g64 );
and ( g_n126 , g119 , g_n122 );
nand ( g_n127 , g_n126 , g43 );
and ( g_n128 , g_n127 , g_n125 );
and ( g_n129 , g119 , g116 );
nand ( g_n130 , g_n129 , g53 );
and ( g_n131 , g_n123 , g116 );
nand ( g_n132 , g_n131 , g32 );
and ( g_n133 , g_n132 , g_n130 );
and ( g_n134 , g_n133 , g_n128 );
or ( g_n135 , g_n134 , g_n121 );
and ( g_n136 , g_n135 , g_n120 );
not ( g_n137 , g134 );
nand ( g_n138 , g144 , g84 );
nand ( g_n139 , g_n82 , g94 );
and ( g_n140 , g_n139 , g145 );
and ( g_n141 , g_n140 , g_n138 );
nand ( g_n142 , g144 , g74 );
nand ( g_n143 , g_n82 , g104 );
and ( g_n144 , g_n143 , g_n83 );
and ( g_n145 , g_n144 , g_n142 );
or ( g_n146 , g_n145 , g_n141 );
or ( g_n147 , g_n146 , g_n137 );
not ( g_n148 , g137 );
nand ( g_n149 , g144 , g91 );
nand ( g_n150 , g_n82 , g101 );
and ( g_n151 , g_n150 , g145 );
and ( g_n152 , g_n151 , g_n149 );
nand ( g_n153 , g144 , g81 );
nand ( g_n154 , g_n82 , g111 );
and ( g_n155 , g_n154 , g_n83 );
and ( g_n156 , g_n155 , g_n153 );
or ( g_n157 , g_n156 , g_n152 );
or ( g_n158 , g_n157 , g_n148 );
and ( g_n159 , g_n158 , g_n147 );
and ( g_n160 , g_n159 , g_n136 );
or ( g_n161 , g_n160 , g_n109 );
and ( g_n162 , g_n106 , g_n94 );
not ( g_n163 , g_n162 );
and ( g_n164 , g_n163 , g7 );
not ( g_n165 , g132 );
nand ( g_n166 , g_n129 , g54 );
nand ( g_n167 , g_n124 , g65 );
and ( g_n168 , g_n167 , g_n166 );
nand ( g_n169 , g_n126 , g44 );
nand ( g_n170 , g_n131 , g33 );
and ( g_n171 , g_n170 , g_n169 );
and ( g_n172 , g_n171 , g_n168 );
or ( g_n173 , g_n172 , g_n165 );
not ( g_n174 , g131 );
nor ( g_n175 , g_n122 , g55 );
or ( g_n176 , g_n175 , g_n123 );
nand ( g_n177 , g_n131 , g34 );
nand ( g_n178 , g_n122 , g66 );
and ( g_n179 , g_n178 , g_n177 );
and ( g_n180 , g_n179 , g_n176 );
or ( g_n181 , g_n180 , g_n174 );
nand ( g_n182 , g_n181 , g_n173 );
nand ( g_n183 , g_n182 , g_n164 );
not ( g_n184 , g_n129 );
nor ( g_n185 , g_n184 , g56 );
not ( g_n186 , g_n131 );
nor ( g_n187 , g_n186 , g35 );
or ( g_n188 , g_n187 , g_n185 );
not ( g_n189 , g_n124 );
nor ( g_n190 , g_n189 , g67 );
not ( g_n191 , g_n126 );
nor ( g_n192 , g_n191 , g45 );
or ( g_n193 , g_n192 , g_n190 );
or ( g_n194 , g_n193 , g_n188 );
nand ( g_n195 , g_n163 , g130 );
nand ( g_n196 , g_n162 , g141 );
and ( g_n197 , g_n196 , g_n195 );
or ( g_n198 , g_n197 , g_n194 );
nor ( g_n199 , g_n191 , g46 );
nor ( g_n200 , g_n186 , g36 );
or ( g_n201 , g_n200 , g_n199 );
nor ( g_n202 , g_n189 , g68 );
nor ( g_n203 , g_n184 , g57 );
or ( g_n204 , g_n203 , g_n202 );
or ( g_n205 , g_n204 , g_n201 );
nand ( g_n206 , g_n163 , g129 );
nand ( g_n207 , g_n162 , g140 );
and ( g_n208 , g_n207 , g_n206 );
or ( g_n209 , g_n208 , g_n205 );
nand ( g_n210 , g_n209 , g_n198 );
nand ( g_n211 , g_n210 , g7 );
nor ( g_n212 , g_n189 , g62 );
nor ( g_n213 , g_n186 , g30 );
or ( g_n214 , g_n213 , g_n212 );
nor ( g_n215 , g_n191 , g41 );
nor ( g_n216 , g_n184 , g51 );
or ( g_n217 , g_n216 , g_n215 );
or ( g_n218 , g_n217 , g_n214 );
not ( g_n219 , g125 );
nor ( g_n220 , g_n189 , g71 );
nor ( g_n221 , g_n186 , g39 );
or ( g_n222 , g_n221 , g_n220 );
nor ( g_n223 , g_n184 , g60 );
nor ( g_n224 , g_n191 , g49 );
or ( g_n225 , g_n224 , g_n223 );
or ( g_n226 , g_n225 , g_n222 );
nor ( g_n227 , g_n226 , g_n219 );
nor ( g_n228 , g_n227 , g124 );
and ( g_n229 , g_n228 , g_n163 );
or ( g_n230 , g_n226 , g_n148 );
and ( g_n231 , g_n230 , g_n110 );
and ( g_n232 , g_n231 , g_n162 );
or ( g_n233 , g_n232 , g_n229 );
and ( g_n234 , g_n233 , g_n218 );
or ( g_n235 , g_n162 , g_n219 );
or ( g_n236 , g_n163 , g_n148 );
and ( g_n237 , g_n236 , g_n226 );
and ( g_n238 , g_n237 , g_n235 );
nand ( g_n239 , g_n126 , g48 );
nand ( g_n240 , g_n129 , g59 );
and ( g_n241 , g_n240 , g_n239 );
nand ( g_n242 , g_n131 , g38 );
nand ( g_n243 , g_n124 , g70 );
and ( g_n244 , g_n243 , g_n242 );
and ( g_n245 , g_n244 , g_n241 );
nand ( g_n246 , g_n163 , g127 );
nand ( g_n247 , g_n162 , g138 );
and ( g_n248 , g_n247 , g_n246 );
and ( g_n249 , g_n248 , g_n245 );
or ( g_n250 , g_n249 , g_n238 );
or ( g_n251 , g_n250 , g_n234 );
nor ( g_n252 , g_n186 , g37 );
nor ( g_n253 , g_n191 , g47 );
or ( g_n254 , g_n253 , g_n252 );
nor ( g_n255 , g_n189 , g69 );
nor ( g_n256 , g_n184 , g58 );
or ( g_n257 , g_n256 , g_n255 );
or ( g_n258 , g_n257 , g_n254 );
nand ( g_n259 , g_n163 , g128 );
nand ( g_n260 , g_n162 , g139 );
and ( g_n261 , g_n260 , g_n259 );
or ( g_n262 , g_n261 , g_n258 );
or ( g_n263 , g_n248 , g_n245 );
and ( g_n264 , g_n263 , g_n262 );
and ( g_n265 , g_n264 , g_n251 );
and ( g_n266 , g_n261 , g_n258 );
and ( g_n267 , g_n205 , g7 );
and ( g_n268 , g_n267 , g_n208 );
or ( g_n269 , g_n268 , g_n266 );
or ( g_n270 , g_n269 , g_n265 );
and ( g_n271 , g_n270 , g_n211 );
and ( g_n272 , g_n194 , g7 );
and ( g_n273 , g_n272 , g_n197 );
or ( g_n274 , g_n273 , g_n271 );
and ( g_n275 , g_n274 , g_n183 );
and ( g_n276 , g_n172 , g_n165 );
and ( g_n277 , g_n180 , g_n174 );
or ( g_n278 , g_n277 , g_n276 );
and ( g_n279 , g_n278 , g_n173 );
and ( g_n280 , g_n279 , g_n164 );
or ( g_n281 , g_n280 , g_n275 );
and ( g_n282 , g_n281 , g_n161 );
or ( g_n283 , g_n120 , g_n109 );
and ( g_n284 , g_n146 , g_n137 );
and ( g_n285 , g_n134 , g_n121 );
or ( g_n286 , g_n285 , g_n284 );
and ( g_n287 , g_n286 , g_n147 );
and ( g_n288 , g_n287 , g_n283 );
and ( g_n289 , g_n157 , g_n148 );
and ( g_n290 , g_n119 , g_n110 );
or ( g_n291 , g_n290 , g_n289 );
or ( g_n292 , g_n291 , g_n288 );
and ( g_n293 , g_n158 , g_n108 );
and ( g_n294 , g_n293 , g_n292 );
endmodule
