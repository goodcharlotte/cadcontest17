module G ( 
    g7 , g29 , g30 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g41 , g43 , g44 ,
    g45 , g46 , g47 , g48 , g49 , g51 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 ,
    g62 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 ,
    g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 ,
    g111 , g112 , g116 , g119 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 ,
    g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 ,
    g217  );
  input  g7 , g29 , g30 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g41 , g43 ,
    g44 , g45 , g46 , g47 , g48 , g49 , g51 , g53 , g54 , g55 , g56 , g57 , g58 , g59 ,
    g60 , g62 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 ,
    g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 ,
    g109 , g111 , g112 , g116 , g119 , g124 , g125 , g126 , g127 , g128 , g129 , g130 ,
    g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 ;
  output g217 ;
  wire n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 ,
    n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 ,
    n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 ,
    n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 ,
    n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 ,
    n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 ,
    n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 ,
    n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 ,
    n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 ,
    n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 ,
    n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 ,
    n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 ,
    n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 ,
    n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 ,
    n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 ,
    n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 ,
    n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 ,
    n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 ;
  and  ( n80 , g145 , g88 );
  not  ( n81 , n80 );
  not  ( n82 , g144 );
  not  ( n83 , g145 );
  and  ( n84 , n83 , g78 );
  nor  ( n85 , n84 , n82 );
  and  ( n86 , n85 , n81 );
  and  ( n87 , g145 , g98 );
  not  ( n88 , n87 );
  and  ( n89 , n83 , g108 );
  nor  ( n90 , n89 , g144 );
  and  ( n91 , n90 , n88 );
  nor  ( n92 , n91 , n86 );
  not  ( n93 , n92 );
  and  ( n94 , n93 , g29 );
  nor  ( n95 , n83 , g89 );
  not  ( n96 , n95 );
  nor  ( n97 , g145 , g79 );
  nor  ( n98 , n97 , n82 );
  and  ( n99 , n98 , n96 );
  nor  ( n100 , n83 , g99 );
  not  ( n101 , n100 );
  nor  ( n102 , g145 , g109 );
  nor  ( n103 , n102 , g144 );
  and  ( n104 , n103 , n101 );
  nor  ( n105 , n104 , n99 );
  nor  ( n106 , n105 , g126 );
  not  ( n107 , n106 );
  and  ( n108 , n107 , n94 );
  not  ( n109 , n108 );
  not  ( n110 , g135 );
  nand  ( n111 , g144 , g92 );
  nand  ( n112 , n82 , g102 );
  and  ( n113 , n112 , g145 );
  and  ( n114 , n113 , n111 );
  nand  ( n115 , g144 , g82 );
  nand  ( n116 , n82 , g112 );
  and  ( n117 , n116 , n83 );
  and  ( n118 , n117 , n115 );
  or  ( n119 , n118 , n114 );
  or  ( n120 , n119 , n110 );
  not  ( n121 , g133 );
  not  ( n122 , g116 );
  not  ( n123 , g119 );
  and  ( n124 , n123 , n122 );
  nand  ( n125 , n124 , g64 );
  and  ( n126 , g119 , n122 );
  nand  ( n127 , n126 , g43 );
  and  ( n128 , n127 , n125 );
  and  ( n129 , g119 , g116 );
  nand  ( n130 , n129 , g53 );
  and  ( n131 , n123 , g116 );
  nand  ( n132 , n131 , g32 );
  and  ( n133 , n132 , n130 );
  and  ( n134 , n133 , n128 );
  or  ( n135 , n134 , n121 );
  and  ( n136 , n135 , n120 );
  not  ( n137 , g134 );
  nand  ( n138 , g144 , g84 );
  nand  ( n139 , n82 , g94 );
  and  ( n140 , n139 , g145 );
  and  ( n141 , n140 , n138 );
  nand  ( n142 , g144 , g74 );
  nand  ( n143 , n82 , g104 );
  and  ( n144 , n143 , n83 );
  and  ( n145 , n144 , n142 );
  or  ( n146 , n145 , n141 );
  or  ( n147 , n146 , n137 );
  not  ( n148 , g137 );
  nand  ( n149 , g144 , g91 );
  nand  ( n150 , n82 , g101 );
  and  ( n151 , n150 , g145 );
  and  ( n152 , n151 , n149 );
  nand  ( n153 , g144 , g81 );
  nand  ( n154 , n82 , g111 );
  and  ( n155 , n154 , n83 );
  and  ( n156 , n155 , n153 );
  or  ( n157 , n156 , n152 );
  or  ( n158 , n157 , n148 );
  and  ( n159 , n158 , n147 );
  and  ( n160 , n159 , n136 );
  or  ( n161 , n160 , n109 );
  and  ( n162 , n106 , n94 );
  not  ( n163 , n162 );
  and  ( n164 , n163 , g7 );
  not  ( n165 , g132 );
  nand  ( n166 , n129 , g54 );
  nand  ( n167 , n124 , g65 );
  and  ( n168 , n167 , n166 );
  nand  ( n169 , n126 , g44 );
  nand  ( n170 , n131 , g33 );
  and  ( n171 , n170 , n169 );
  and  ( n172 , n171 , n168 );
  or  ( n173 , n172 , n165 );
  not  ( n174 , g131 );
  nor  ( n175 , n122 , g55 );
  or  ( n176 , n175 , n123 );
  nand  ( n177 , n131 , g34 );
  nand  ( n178 , n122 , g66 );
  and  ( n179 , n178 , n177 );
  and  ( n180 , n179 , n176 );
  or  ( n181 , n180 , n174 );
  nand  ( n182 , n181 , n173 );
  nand  ( n183 , n182 , n164 );
  not  ( n184 , n129 );
  nor  ( n185 , n184 , g56 );
  not  ( n186 , n131 );
  nor  ( n187 , n186 , g35 );
  or  ( n188 , n187 , n185 );
  not  ( n189 , n124 );
  nor  ( n190 , n189 , g67 );
  not  ( n191 , n126 );
  nor  ( n192 , n191 , g45 );
  or  ( n193 , n192 , n190 );
  or  ( n194 , n193 , n188 );
  nand  ( n195 , n163 , g130 );
  nand  ( n196 , n162 , g141 );
  and  ( n197 , n196 , n195 );
  or  ( n198 , n197 , n194 );
  nor  ( n199 , n191 , g46 );
  nor  ( n200 , n186 , g36 );
  or  ( n201 , n200 , n199 );
  nor  ( n202 , n189 , g68 );
  nor  ( n203 , n184 , g57 );
  or  ( n204 , n203 , n202 );
  or  ( n205 , n204 , n201 );
  nand  ( n206 , n163 , g129 );
  nand  ( n207 , n162 , g140 );
  and  ( n208 , n207 , n206 );
  or  ( n209 , n208 , n205 );
  nand  ( n210 , n209 , n198 );
  nand  ( n211 , n210 , g7 );
  nor  ( n212 , n189 , g62 );
  nor  ( n213 , n186 , g30 );
  or  ( n214 , n213 , n212 );
  nor  ( n215 , n191 , g41 );
  nor  ( n216 , n184 , g51 );
  or  ( n217 , n216 , n215 );
  or  ( n218 , n217 , n214 );
  not  ( n219 , g125 );
  nor  ( n220 , n189 , g71 );
  nor  ( n221 , n186 , g39 );
  or  ( n222 , n221 , n220 );
  nor  ( n223 , n184 , g60 );
  nor  ( n224 , n191 , g49 );
  or  ( n225 , n224 , n223 );
  or  ( n226 , n225 , n222 );
  nor  ( n227 , n226 , n219 );
  nor  ( n228 , n227 , g124 );
  and  ( n229 , n228 , n163 );
  or  ( n230 , n226 , n148 );
  and  ( n231 , n230 , n110 );
  and  ( n232 , n231 , n162 );
  or  ( n233 , n232 , n229 );
  and  ( n234 , n233 , n218 );
  or  ( n235 , n162 , n219 );
  or  ( n236 , n163 , n148 );
  and  ( n237 , n236 , n226 );
  and  ( n238 , n237 , n235 );
  nand  ( n239 , n126 , g48 );
  nand  ( n240 , n129 , g59 );
  and  ( n241 , n240 , n239 );
  nand  ( n242 , n131 , g38 );
  nand  ( n243 , n124 , g70 );
  and  ( n244 , n243 , n242 );
  and  ( n245 , n244 , n241 );
  nand  ( n246 , n163 , g127 );
  nand  ( n247 , n162 , g138 );
  and  ( n248 , n247 , n246 );
  and  ( n249 , n248 , n245 );
  or  ( n250 , n249 , n238 );
  or  ( n251 , n250 , n234 );
  nor  ( n252 , n186 , g37 );
  nor  ( n253 , n191 , g47 );
  or  ( n254 , n253 , n252 );
  nor  ( n255 , n189 , g69 );
  nor  ( n256 , n184 , g58 );
  or  ( n257 , n256 , n255 );
  or  ( n258 , n257 , n254 );
  nand  ( n259 , n163 , g128 );
  nand  ( n260 , n162 , g139 );
  and  ( n261 , n260 , n259 );
  or  ( n262 , n261 , n258 );
  or  ( n263 , n248 , n245 );
  and  ( n264 , n263 , n262 );
  and  ( n265 , n264 , n251 );
  and  ( n266 , n261 , n258 );
  and  ( n267 , n205 , g7 );
  and  ( n268 , n267 , n208 );
  or  ( n269 , n268 , n266 );
  or  ( n270 , n269 , n265 );
  and  ( n271 , n270 , n211 );
  and  ( n272 , n194 , g7 );
  and  ( n273 , n272 , n197 );
  or  ( n274 , n273 , n271 );
  and  ( n275 , n274 , n183 );
  and  ( n276 , n172 , n165 );
  and  ( n277 , n180 , n174 );
  or  ( n278 , n277 , n276 );
  and  ( n279 , n278 , n173 );
  and  ( n280 , n279 , n164 );
  or  ( n281 , n280 , n275 );
  and  ( n282 , n281 , n161 );
  or  ( n283 , n120 , n109 );
  and  ( n284 , n146 , n137 );
  and  ( n285 , n134 , n121 );
  or  ( n286 , n285 , n284 );
  and  ( n287 , n286 , n147 );
  and  ( n288 , n287 , n283 );
  and  ( n289 , n157 , n148 );
  and  ( n290 , n119 , n110 );
  or  ( n291 , n290 , n289 );
  or  ( n292 , n291 , n288 );
  and  ( n293 , n158 , n108 );
  and  ( n294 , n293 , n292 );
  or  ( g217 , n294 , n282 );
endmodule


