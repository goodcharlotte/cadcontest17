module  patch (g7 , g29 , g30 , g35 , g41 , g45 , g51 , g56 , g62 , g67 , g116 , g119 , g124 , g125 , g129 , g131 , g132 , g133 , g134 , g135 , g137 , g140 , n89 , n91 , n93 , n94 , n102 , n106 , n114 , n117 , n124 , n142 , n149 , n163 , n171 , n177 , n184 , n196 , n211 , n216 , t_0 );
input g7 , g29 , g30 , g35 , g41 , g45 , g51 , g56 , g62 , g67 , g116 , g119 , g124 , g125 , g129 , g131 , g132 , g133 , g134 , g135 , g137 , g140 , n89 , n91 , n93 , n94 , n102 , n106 , n114 , n117 , n124 , n142 , n149 , n163 , n171 , n177 , n184 , n196 , n211 , n216 ;
output t_0 ;
wire n81 , n82 , n83 , n84 , n85 , n86 , n87 , n104 , n107 , n108 , n109 , n118 , n119 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n143 , n144 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n164 , n172 , n178 , n179 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n197 , n198 , n199 , n200 , n201 , n202 , n212 , n213 , n214 , n215 , n217 , INV_g116 , INV_g119 , INV_g129 , INV_g131 , INV_g132 , INV_g135 , INV_g137 , INV_g140 , INV_n89 , INV_n91 , INV_n93 , INV_n94 , INV_n102 , INV_n106 , INV_n142 , INV_n171 , INV_n177 , INV_n211 , INV_n216 ;
and ( t_0 , n217 , n191 , n137 , n108 );
not ( n81 , INV_g116 );
not ( n82 , INV_g119 );
nor ( n83 , n82 , n81 , g56 );
nor ( n84 , n82 , INV_g116 , g45 );
nor ( n85 , INV_g119 , n81 , g35 );
nor ( n86 , INV_g119 , INV_g116 , g67 );
nor ( n87 , n86 , n85 , n84 , n83 , n80 );
not ( n104 , INV_n102 );
not ( n107 , INV_n106 );
nand ( n108 , n107 , n87 );
or ( n109 , n107 , n87 );
not ( n118 , n117 );
nand ( n119 , n118 , n114 );
and ( n125 , n124 , g125 );
nor ( n126 , n125 , g124 );
or ( n127 , n126 , INV_n102 );
not ( n128 , INV_g135 );
nand ( n129 , n124 , INV_g137 );
and ( n130 , n129 , n128 );
or ( n131 , n130 , n104 );
nor ( n132 , INV_g119 , INV_g116 , g62 );
nor ( n133 , INV_g119 , n81 , g30 );
nor ( n134 , n82 , INV_g116 , g41 );
nor ( n135 , n82 , n81 , g51 );
or ( n136 , n135 , n134 , n133 , n132 );
and ( n137 , n136 , n131 , n127 , n119 , n109 );
not ( n143 , INV_n142 );
nand ( n144 , n143 , INV_g132 );
not ( n150 , n149 );
nand ( n151 , n150 , INV_g131 );
or ( n152 , n143 , INV_g132 );
or ( n153 , n150 , INV_g131 );
and ( n154 , n153 , n152 , n151 , n144 );
or ( n155 , n154 , n80 );
not ( n156 , g134 );
nand ( n164 , n163 , n156 );
or ( n172 , INV_n171 , n128 );
xor ( n178 , INV_n177 , INV_g137 );
and ( n179 , n178 , n172 , n164 );
xor ( n185 , n184 , g133 );
nand ( n186 , INV_n171 , n128 );
or ( n187 , n163 , n156 );
and ( n188 , n187 , n186 , n185 , n179 );
or ( n189 , n188 , n96 );
and ( n190 , n189 , n155 );
or ( n191 , n190 , INV_n102 );
and ( n197 , n104 , INV_g129 );
and ( n198 , INV_n102 , INV_g140 );
nor ( n199 , n198 , n197 );
and ( n200 , n199 , n196 );
nor ( n201 , n199 , n196 );
or ( n202 , n201 , n200 , n80 );
or ( n212 , n118 , n114 );
and ( n213 , n104 , g125 );
and ( n214 , INV_n102 , INV_g137 );
or ( n215 , n214 , n213 , n124 );
and ( n217 , INV_n216 , n215 , n212 , INV_n211 , n202 );
not ( INV_g116 , g116 );
not ( INV_g119 , g119 );
not ( INV_g129 , g129 );
not ( INV_g131 , g131 );
not ( INV_g132 , g132 );
not ( INV_g135 , g135 );
not ( INV_g137 , g137 );
not ( INV_g140 , g140 );
not ( INV_n89 , n89 );
not ( INV_n91 , n91 );
not ( INV_n93 , n93 );
not ( INV_n94 , n94 );
not ( INV_n102 , n102 );
not ( INV_n106 , n106 );
not ( INV_n142 , n142 );
not ( INV_n171 , n171 );
not ( INV_n177 , n177 );
not ( INV_n211 , n211 );
not ( INV_n216 , n216 );
endmodule
