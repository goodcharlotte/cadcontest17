module F ( 
    g7 , g29 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g43 , g44 , g45 , g46 ,
    g47 , g48 , g49 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g64 , g65 , g66 ,
    g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 ,
    g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 ,
    g119 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 ,
    g137 , g138 , g139 , g140 , g141 , g144 , g145 , t_0 ,
    g217  );
  input  g7 , g29 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g43 , g44 , g45 ,
    g46 , g47 , g48 , g49 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g64 , g65 ,
    g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 ,
    g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 ,
    g116 , g119 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 ,
    g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 , t_0 ;
  output g217 ;
  wire n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 ,
    n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 ,
    n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ,
    n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 ,
    n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 ,
    n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 ,
    n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 ,
    n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 ,
    n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 ,
    n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 ,
    n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 ,
    n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 ,
    n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 ,
    n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 ,
    n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 ,
    n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 ,
    n271 , n272 , n273 , n274 , n275 ;
  assign n76 = ~g144 & g145;
  assign n77 = g94 & n76;
  assign n78 = g144 & g145;
  assign n79 = g84 & n78;
  assign n80 = g144 & ~g145;
  assign n81 = g74 & n80;
  assign n82 = ~g144 & ~g145;
  assign n83 = g104 & n82;
  assign n84 = ~n77 & ~n79;
  assign n85 = ~n81 & ~n83;
  assign n86 = n84 & n85;
  assign n87 = g99 & n76;
  assign n88 = g79 & n80;
  assign n89 = g89 & n78;
  assign n90 = g109 & n82;
  assign n91 = ~n87 & ~n88;
  assign n92 = ~n89 & ~n90;
  assign n93 = n91 & n92;
  assign n94 = ~g126 & ~n93;
  assign n95 = g78 & n80;
  assign n96 = g108 & n82;
  assign n97 = g88 & n78;
  assign n98 = g98 & n76;
  assign n99 = g29 & ~n95;
  assign n100 = ~n96 & ~n97;
  assign n101 = ~n98 & n100;
  assign n102 = n99 & n101;
  assign n103 = ~n94 & n102;
  assign n104 = g134 & ~n86;
  assign n105 = n103 & n104;
  assign n106 = g81 & n80;
  assign n107 = g91 & n78;
  assign n108 = g111 & n82;
  assign n109 = g101 & n76;
  assign n110 = ~n106 & ~n107;
  assign n111 = ~n108 & ~n109;
  assign n112 = n110 & n111;
  assign n113 = n103 & ~n112;
  assign n114 = g137 & n113;
  assign n115 = ~g137 & n103;
  assign n116 = ~n113 & n115;
  assign n117 = ~n114 & ~n116;
  assign n118 = ~g134 & n86;
  assign n119 = n103 & n118;
  assign n120 = ~n105 & ~n119;
  assign n121 = n117 & n120;
  assign n122 = n94 & n102;
  assign n123 = g7 & ~n122;
  assign n124 = g34 & ~g119;
  assign n125 = g55 & g119;
  assign n126 = g116 & ~n124;
  assign n127 = ~n125 & n126;
  assign n128 = ~g66 & ~g116;
  assign n129 = ~g119 & n128;
  assign n130 = ~n127 & ~n129;
  assign n131 = ~g131 & ~n130;
  assign n132 = ~g44 & ~g116;
  assign n133 = ~g54 & g116;
  assign n134 = g119 & ~n132;
  assign n135 = ~n133 & n134;
  assign n136 = ~g65 & ~g116;
  assign n137 = ~g33 & g116;
  assign n138 = ~g119 & ~n136;
  assign n139 = ~n137 & n138;
  assign n140 = ~n135 & ~n139;
  assign n141 = g132 & ~n140;
  assign n142 = n123 & n141;
  assign n143 = n123 & n131;
  assign n144 = ~n142 & n143;
  assign n145 = ~g132 & n140;
  assign n146 = n123 & n145;
  assign n147 = g140 & n122;
  assign n148 = g129 & ~n122;
  assign n149 = ~g46 & ~g116;
  assign n150 = ~g57 & g116;
  assign n151 = g119 & ~n149;
  assign n152 = ~n150 & n151;
  assign n153 = ~g68 & ~g116;
  assign n154 = ~g36 & g116;
  assign n155 = ~g119 & ~n153;
  assign n156 = ~n154 & n155;
  assign n157 = ~n152 & ~n156;
  assign n158 = g7 & ~n157;
  assign n159 = ~g37 & ~g119;
  assign n160 = ~g58 & g119;
  assign n161 = g116 & ~n159;
  assign n162 = ~n160 & n161;
  assign n163 = ~g69 & ~g119;
  assign n164 = ~g47 & g119;
  assign n165 = ~g116 & ~n163;
  assign n166 = ~n164 & n165;
  assign n167 = ~n162 & ~n166;
  assign n168 = g128 & ~n122;
  assign n169 = g139 & n122;
  assign n170 = ~n168 & ~n169;
  assign n171 = ~n167 & ~n170;
  assign n172 = n167 & n170;
  assign n173 = ~g48 & ~g116;
  assign n174 = ~g59 & g116;
  assign n175 = g119 & ~n173;
  assign n176 = ~n174 & n175;
  assign n177 = ~g70 & ~g116;
  assign n178 = ~g38 & g116;
  assign n179 = ~g119 & ~n177;
  assign n180 = ~n178 & n179;
  assign n181 = ~n176 & ~n180;
  assign n182 = g127 & ~n122;
  assign n183 = g138 & n122;
  assign n184 = ~n182 & ~n183;
  assign n185 = ~n181 & ~n184;
  assign n186 = n181 & n184;
  assign n187 = ~g49 & ~g116;
  assign n188 = ~g60 & g116;
  assign n189 = g119 & ~n187;
  assign n190 = ~n188 & n189;
  assign n191 = ~g71 & ~g116;
  assign n192 = ~g39 & g116;
  assign n193 = ~g119 & ~n191;
  assign n194 = ~n192 & n193;
  assign n195 = ~n190 & ~n194;
  assign n196 = ~t_0 & ~n195;
  assign n197 = t_0 & n195;
  assign n198 = g125 & ~n122;
  assign n199 = g137 & n122;
  assign n200 = ~n198 & ~n199;
  assign n201 = ~n197 & ~n200;
  assign n202 = ~n196 & ~n201;
  assign n203 = ~n186 & ~n202;
  assign n204 = ~n185 & ~n203;
  assign n205 = ~n172 & ~n204;
  assign n206 = ~n171 & ~n205;
  assign n207 = n158 & ~n206;
  assign n208 = g7 & ~n147;
  assign n209 = ~n148 & n208;
  assign n210 = ~n207 & n209;
  assign n211 = ~g45 & ~g116;
  assign n212 = ~g56 & g116;
  assign n213 = g119 & ~n211;
  assign n214 = ~n212 & n213;
  assign n215 = ~g67 & ~g116;
  assign n216 = ~g35 & g116;
  assign n217 = ~g119 & ~n215;
  assign n218 = ~n216 & n217;
  assign n219 = ~n214 & ~n218;
  assign n220 = g7 & ~n219;
  assign n221 = g141 & n122;
  assign n222 = g130 & ~n122;
  assign n223 = g7 & ~n221;
  assign n224 = ~n222 & n223;
  assign n225 = ~n220 & n224;
  assign n226 = ~n158 & n206;
  assign n227 = ~n225 & ~n226;
  assign n228 = ~n210 & n227;
  assign n229 = g131 & n130;
  assign n230 = ~n131 & ~n229;
  assign n231 = n123 & ~n230;
  assign n232 = n220 & ~n224;
  assign n233 = ~n142 & ~n146;
  assign n234 = ~n231 & n233;
  assign n235 = ~n232 & n234;
  assign n236 = ~n228 & n235;
  assign n237 = ~n144 & ~n146;
  assign n238 = ~n236 & n237;
  assign n239 = ~g43 & ~g116;
  assign n240 = ~g53 & g116;
  assign n241 = g119 & ~n239;
  assign n242 = ~n240 & n241;
  assign n243 = ~g64 & ~g116;
  assign n244 = ~g32 & g116;
  assign n245 = ~g119 & ~n243;
  assign n246 = ~n244 & n245;
  assign n247 = ~n242 & ~n246;
  assign n248 = ~g133 & n247;
  assign n249 = n103 & n248;
  assign n250 = g102 & n76;
  assign n251 = g92 & n78;
  assign n252 = g82 & n80;
  assign n253 = g112 & n82;
  assign n254 = ~n250 & ~n251;
  assign n255 = ~n252 & ~n253;
  assign n256 = n254 & n255;
  assign n257 = n103 & ~n256;
  assign n258 = g135 & n257;
  assign n259 = ~g135 & n103;
  assign n260 = ~n257 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = g133 & ~n247;
  assign n263 = n103 & n262;
  assign n264 = ~n249 & ~n263;
  assign n265 = n261 & n264;
  assign n266 = n121 & n265;
  assign n267 = ~n238 & n266;
  assign n268 = ~n114 & n260;
  assign n269 = n249 & n261;
  assign n270 = n121 & n269;
  assign n271 = n117 & n119;
  assign n272 = n261 & n271;
  assign n273 = ~n116 & ~n268;
  assign n274 = ~n270 & n273;
  assign n275 = ~n272 & n274;
  assign g217 = n267 | ~n275;
endmodule


