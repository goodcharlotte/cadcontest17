module F ( g7 , g29 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 , g119 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 , t_0 , g217 );
input g7 , g29 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 , g119 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 , t_0 ;
output g217 ;
wire n8 , n30 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n75 , n79 , n80 , n82 , n83 , n85 , n89 , n90 , n92 , n93 , n95 , n99 , n100 , n102 , n103 , n105 , n109 , n110 , n112 , n113 , n117 , n120 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , n145 , n146 , n218 , n477 , n373 , n244 , n378 , n400 , n348 , n448 , n494 , n588 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n318 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n374 , n375 , n376 , n377 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 ;
buf ( g217 , n218 );
buf ( n8 , g7 );
buf ( n30 , g29 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n75 , g74 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n85 , g84 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n95 , g94 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n105 , g104 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n117 , g116 );
buf ( n120 , g119 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n218 , n588 );
not ( n477 , n476 );
nor ( n373 , n366 , n372 );
nand ( n244 , n237 , n243 );
nand ( n378 , n376 , n377 , n371 );
nand ( n400 , n395 , n399 );
not ( n348 , n347 );
nand ( n448 , n439 , n447 );
nand ( n494 , n490 , n492 , n493 );
nor ( n588 , n584 , n587 );
not ( n229 , n49 );
not ( n230 , n117 );
nand ( n231 , n230 , n120 );
not ( n232 , n231 );
not ( n233 , n232 );
or ( n234 , n229 , n233 );
nand ( n235 , n120 , n60 , n117 );
nand ( n236 , n234 , n235 );
not ( n237 , n236 );
not ( n238 , n120 );
and ( n239 , n117 , n39 );
not ( n240 , n117 );
and ( n241 , n240 , n71 );
or ( n242 , n239 , n241 );
nand ( n243 , n238 , n242 );
not ( n245 , n244 );
not ( n246 , n146 );
not ( n247 , n246 );
not ( n248 , n110 );
nor ( n249 , n248 , n145 );
not ( n250 , n249 );
or ( n251 , n247 , n250 );
nand ( n252 , n146 , n90 , n145 );
nand ( n253 , n251 , n252 );
not ( n254 , n145 );
nand ( n255 , n254 , n146 , n100 );
not ( n256 , n146 );
nand ( n257 , n256 , n80 , n145 );
nand ( n258 , n255 , n257 );
nor ( n259 , n253 , n258 );
not ( n260 , n259 );
not ( n261 , n146 );
nand ( n262 , n261 , n79 , n145 );
not ( n263 , n145 );
nand ( n264 , n263 , n146 , n99 );
nand ( n265 , n262 , n264 );
not ( n266 , n146 );
not ( n267 , n109 );
nor ( n268 , n267 , n145 );
nand ( n269 , n266 , n268 );
nand ( n270 , n146 , n89 , n145 );
nand ( n271 , n269 , n270 );
nor ( n272 , n265 , n271 );
not ( n273 , n127 );
and ( n274 , n260 , n272 , n273 , n30 );
buf ( n275 , n274 );
and ( n276 , n275 , n139 );
not ( n277 , n275 );
and ( n278 , n277 , n128 );
nor ( n279 , n276 , n278 );
not ( n280 , n279 );
or ( n281 , n245 , n280 );
or ( n282 , n244 , n279 );
nand ( n283 , n281 , n282 );
and ( n284 , n275 , n138 );
not ( n285 , n275 );
and ( n286 , n285 , n126 );
nor ( n287 , n284 , n286 );
nand ( n288 , n61 , n117 );
and ( n289 , n120 , n288 );
not ( n290 , n120 );
not ( n291 , n117 );
nand ( n292 , n291 , n72 );
and ( n293 , n290 , n292 );
or ( n294 , n289 , n293 );
not ( n295 , n120 );
nand ( n296 , n295 , n40 , n117 );
not ( n297 , n231 );
nand ( n298 , n50 , n297 );
nand ( n299 , n294 , n296 , n298 );
not ( n300 , n299 );
not ( n301 , n300 );
not ( n302 , n301 );
not ( n303 , n302 );
not ( n304 , n303 );
nand ( n305 , n283 , n287 , n304 );
not ( n306 , n243 );
nor ( n307 , n236 , n306 );
nand ( n308 , n307 , n279 );
not ( n318 , n117 );
not ( n322 , n136 );
not ( n323 , n303 );
not ( n324 , n287 );
or ( n325 , n323 , n324 );
or ( n326 , n303 , n287 );
nand ( n327 , n325 , n326 );
nand ( n328 , t_0 , n327 , n283 );
nand ( n329 , n305 , n308 , n328 );
nor ( n330 , n259 , n127 );
and ( n331 , n330 , n272 , n30 );
not ( n332 , n331 );
not ( n333 , n132 );
nand ( n334 , n332 , n333 , n8 );
not ( n335 , n334 );
not ( n336 , n335 );
not ( n337 , n275 );
nand ( n338 , n120 , n318 );
not ( n339 , n338 );
not ( n340 , n339 );
nand ( n341 , n120 , n56 , n117 );
not ( n342 , n120 );
nand ( n343 , n342 , n35 , n117 );
not ( n344 , n120 );
nand ( n345 , n344 , n67 , n318 );
nand ( n346 , n340 , n341 , n343 , n345 );
not ( n347 , n346 );
nand ( n349 , n337 , n8 , n348 );
not ( n350 , n349 );
not ( n351 , n350 );
or ( n352 , n336 , n351 );
nand ( n353 , n334 , n349 );
nand ( n354 , n352 , n353 );
not ( n355 , n275 );
or ( n356 , n140 , n355 );
not ( n357 , n129 );
not ( n358 , n275 );
nand ( n359 , n357 , n358 );
nand ( n360 , n356 , n359 );
nand ( n361 , n59 , n117 );
and ( n362 , n120 , n361 );
not ( n363 , n120 );
nand ( n364 , n38 , n117 );
and ( n365 , n363 , n364 );
nor ( n366 , n362 , n365 );
not ( n367 , n48 );
not ( n368 , n297 );
or ( n369 , n367 , n368 );
not ( n370 , n120 );
nand ( n371 , n370 , n70 , n318 );
nand ( n372 , n369 , n371 );
and ( n374 , n360 , n373 );
not ( n375 , n360 );
not ( n376 , n366 );
nand ( n377 , n48 , n339 );
and ( n379 , n375 , n378 );
nor ( n380 , n374 , n379 );
not ( n381 , n131 );
nor ( n382 , n381 , n331 );
not ( n383 , n142 );
not ( n384 , n331 );
or ( n385 , n383 , n384 );
nand ( n386 , n385 , n8 );
nor ( n387 , n382 , n386 );
not ( n388 , n46 );
not ( n389 , n338 );
not ( n390 , n389 );
or ( n391 , n388 , n390 );
not ( n392 , n120 );
nand ( n393 , n392 , n36 , n117 );
nand ( n394 , n391 , n393 );
not ( n395 , n394 );
nand ( n396 , n120 , n57 , n117 );
not ( n397 , n120 );
nand ( n398 , n397 , n68 , n318 );
and ( n399 , n396 , n398 );
nand ( n401 , n8 , n400 );
not ( n402 , n401 );
and ( n403 , n387 , n402 );
not ( n404 , n387 );
and ( n405 , n404 , n401 );
nor ( n406 , n403 , n405 );
not ( n407 , n406 );
nand ( n408 , n354 , n380 , n407 );
not ( n409 , n141 );
not ( n410 , n331 );
or ( n411 , n409 , n410 );
nand ( n412 , n411 , n8 );
not ( n413 , n130 );
nor ( n414 , n413 , n331 );
nor ( n415 , n412 , n414 );
and ( n416 , n120 , n58 , n117 );
not ( n417 , n69 );
nor ( n418 , n417 , n120 , n117 );
nor ( n419 , n416 , n418 );
nand ( n420 , n37 , n117 );
nor ( n421 , n120 , n420 );
not ( n422 , n421 );
nand ( n423 , n47 , n339 );
nand ( n424 , n419 , n422 , n423 );
nand ( n425 , n8 , n424 );
and ( n426 , n415 , n425 );
not ( n427 , n415 );
not ( n428 , n425 );
and ( n429 , n427 , n428 );
nor ( n430 , n426 , n429 );
not ( n431 , n331 );
not ( n432 , n133 );
nand ( n433 , n431 , n432 , n8 );
not ( n434 , n433 );
not ( n435 , n275 );
and ( n436 , n45 , n232 );
nand ( n437 , n34 , n117 );
nor ( n438 , n120 , n437 );
nor ( n439 , n436 , n438 );
nand ( n440 , n55 , n117 );
not ( n441 , n440 );
and ( n442 , n120 , n441 );
not ( n443 , n120 );
not ( n444 , n66 );
nor ( n445 , n444 , n117 );
and ( n446 , n443 , n445 );
nor ( n447 , n442 , n446 );
nand ( n449 , n435 , n8 , n448 );
xor ( n450 , n434 , n449 );
nand ( n451 , n430 , n450 );
nor ( n452 , n408 , n451 );
and ( n453 , n329 , n452 );
nand ( n454 , n407 , n430 );
nand ( n455 , n373 , n360 );
nand ( n456 , n354 , n450 );
nor ( n457 , n454 , n455 , n456 );
nor ( n458 , n453 , n457 );
and ( n459 , n450 , n335 , n349 );
and ( n460 , n434 , n449 );
nor ( n461 , n459 , n460 );
not ( n462 , n461 );
nand ( n463 , n415 , n450 );
not ( n464 , n406 );
nand ( n465 , n464 , n354 , n425 );
nor ( n466 , n463 , n465 );
buf ( n467 , n387 );
nand ( n468 , n354 , n467 );
nand ( n469 , n401 , n450 );
nor ( n470 , n468 , n469 );
nor ( n471 , n462 , n466 , n470 );
nand ( n472 , n458 , n471 );
not ( n473 , n134 );
not ( n474 , n330 );
nor ( n475 , n265 , n271 );
not ( n476 , n475 );
nand ( n478 , n474 , n477 , n30 );
not ( n479 , n478 );
not ( n480 , n275 );
and ( n481 , n473 , n479 , n480 );
not ( n482 , n481 );
nand ( n483 , n54 , n117 );
not ( n484 , n483 );
and ( n485 , n120 , n484 );
not ( n486 , n120 );
not ( n487 , n65 );
nor ( n488 , n487 , n117 );
and ( n489 , n486 , n488 );
nor ( n490 , n485 , n489 );
not ( n491 , n120 );
nand ( n492 , n491 , n33 , n117 );
nand ( n493 , n44 , n339 );
and ( n495 , n494 , n479 , n480 );
not ( n496 , n495 );
or ( n497 , n482 , n496 );
or ( n498 , n481 , n495 );
nand ( n499 , n497 , n498 );
not ( n500 , n135 );
and ( n501 , n500 , n479 , n355 );
not ( n502 , n275 );
not ( n503 , n95 );
not ( n504 , n146 );
nor ( n505 , n504 , n145 );
not ( n506 , n505 );
or ( n507 , n503 , n506 );
nand ( n508 , n145 , n146 );
not ( n509 , n508 );
nand ( n510 , n85 , n509 );
nand ( n511 , n507 , n510 );
not ( n512 , n75 );
not ( n513 , n145 );
nor ( n514 , n513 , n146 );
not ( n515 , n514 );
or ( n516 , n512 , n515 );
nor ( n517 , n145 , n146 );
nand ( n518 , n105 , n517 );
nand ( n519 , n516 , n518 );
nor ( n520 , n511 , n519 );
not ( n521 , n520 );
nand ( n522 , n502 , n521 , n479 );
xor ( n523 , n501 , n522 );
not ( n524 , n275 );
not ( n525 , n138 );
nand ( n526 , n524 , n525 , n479 );
not ( n527 , n526 );
not ( n528 , n527 );
not ( n529 , n275 );
not ( n530 , n92 );
not ( n531 , n530 );
nand ( n532 , n145 , n146 );
not ( n533 , n532 );
and ( n534 , n531 , n533 );
nor ( n535 , n145 , n146 );
and ( n536 , n112 , n535 );
nor ( n537 , n534 , n536 );
not ( n538 , n146 );
nor ( n539 , n538 , n145 );
nand ( n540 , n102 , n539 );
not ( n541 , n145 );
nor ( n542 , n541 , n146 );
nand ( n543 , n82 , n542 );
nand ( n544 , n537 , n540 , n543 );
not ( n545 , n544 );
not ( n546 , n545 );
nand ( n547 , n529 , n546 , n479 );
not ( n548 , n547 );
not ( n549 , n548 );
or ( n550 , n528 , n549 );
nand ( n551 , n526 , n547 );
nand ( n552 , n550 , n551 );
not ( n553 , n275 );
nand ( n554 , n553 , n322 , n479 );
not ( n555 , n554 );
not ( n556 , n555 );
and ( n557 , n103 , n539 );
not ( n558 , n93 );
nor ( n559 , n558 , n532 );
nor ( n560 , n557 , n559 );
and ( n561 , n83 , n542 );
and ( n562 , n113 , n517 );
nor ( n563 , n561 , n562 );
nand ( n564 , n560 , n563 );
and ( n565 , n564 , n479 , n355 );
not ( n566 , n565 );
or ( n567 , n556 , n566 );
or ( n568 , n555 , n565 );
nand ( n569 , n567 , n568 );
and ( n570 , n499 , n523 , n552 , n569 );
not ( n571 , n565 );
nand ( n572 , n552 , n571 , n555 );
and ( n573 , n501 , n522 );
nand ( n574 , n573 , n552 , n569 );
and ( n575 , n572 , n574 );
nand ( n576 , n527 , n547 );
nand ( n577 , n481 , n552 , n523 );
not ( n578 , n577 );
not ( n579 , n569 );
nor ( n580 , n579 , n495 );
nand ( n581 , n578 , n580 );
nand ( n582 , n575 , n576 , n581 );
nor ( n583 , n570 , n582 );
and ( n584 , n472 , n583 );
not ( n585 , n472 );
not ( n586 , n582 );
and ( n587 , n585 , n586 );
endmodule
