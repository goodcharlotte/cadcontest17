module G ( g7 , g29 , g30 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g41 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g51 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g62 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 , g119 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 , g217 );
input g7 , g29 , g30 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g41 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g51 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g62 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g74 , g78 , g79 , g81 , g82 , g84 , g88 , g89 , g91 , g92 , g94 , g98 , g99 , g101 , g102 , g104 , g108 , g109 , g111 , g112 , g116 , g119 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g137 , g138 , g139 , g140 , g141 , g144 , g145 ;
output g217 ;
wire g4676 , g4698 , g4699 , g4701 , g4702 , g4703 , g4704 , g4705 , g4706 , g4707 , g4708 , g4710 , g4712 , g4713 , g4714 , g4715 , g4716 , g4717 , g4718 , g4720 , g4722 , g4723 , g4724 , g4725 , g4726 , g4727 , g4728 , g4729 , g4731 , g4733 , g4734 , g4735 , g4736 , g4737 , g4738 , g4739 , g4740 , g4743 , g4747 , g4748 , g4750 , g4751 , g4753 , g4757 , g4758 , g4760 , g4761 , g4763 , g4767 , g4768 , g4770 , g4771 , g4773 , g4777 , g4778 , g4780 , g4781 , g4785 , g4788 , g4793 , g4794 , g4795 , g4796 , g4797 , g4798 , g4799 , g4800 , g4801 , g4802 , g4803 , g4804 , g4806 , g4807 , g4808 , g4809 , g4810 , g4813 , g4814 , g4886 , g807 , g653 , g589 , g975 , g1199 , g1245 , g732 , g1135 , g457 , g1377 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g466 , g488 , g489 , g495 , g501 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g550 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g607 , g608 , g609 , g610 , g611 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g658 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g685 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g720 , g725 , g726 , g727 , g728 , g729 , g730 , g731 , g739 , g750 , g771 , g790 , g794 , g795 , g796 , g797 , g798 , g799 , g800 , g801 , g802 , g803 , g804 , g805 , g806 , g813 , g822 , g823 , g824 , g825 , g826 , g827 , g828 , g829 , g830 , g831 , g832 , g833 , g834 , g835 , g836 , g837 , g838 , g839 , g840 , g841 , g842 , g843 , g844 , g845 , g846 , g847 , g848 , g849 , g850 , g851 , g852 , g853 , g854 , g855 , g856 , g857 , g858 , g859 , g860 , g861 , g862 , g863 , g869 , g870 , g960 , g961 , g962 , g963 , g964 , g965 , g966 , g967 , g968 , g969 , g970 , g977 , g978 , g979 , g980 , g1005 , g1006 , g1007 , g1008 , g1009 , g1010 , g1011 , g1134 , g1136 , g1137 , g1138 , g1246 , g1247 , g1248 , g1249 , g1250 , g1251 , g1252 , g1253 , g1254 , g1255 , g1256 , g1257 , g1258 , g1259 , g1265 , g1266 , g1267 , g1268 , g1269 , g1270 , g1271 , g1272 , g1273 , g1274 , g1275 , g1276 , g1277 , g1278 , g1279 , g1280 , g1281 , g1282 , g1283 , g1284 , g1285 , g1286 , g1287 , g1288 , g1289 , g1290 , g1291 , g1292 , g1293 , g1294 , g1295 , g1296 , g1297 , g1298 , g1299 , g1300 , g1301 , g1302 , g1303 , g1304 , g1305 , g1306 , g1307 , g1308 , g1309 , g1310 , g1311 , g1312 , g1313 , g1314 , g1315 , g1316 , g1317 , g1318 , g1319 , g1320 , g1321 , g1326 , g1327 , g1328 , g1329 , g1330 , g1331 , g1332 , g1333 , g1334 , g1335 , g1349 , g1359 , g1360 , g1361 , g1362 , g1363 , g1364 , g1365 , g1366 , g1367 , g1368 , g1369 , g1370 , g1371 , g1372 , g1373 , g1374 , g1375 , g1376 ;
buf ( g217 , g4886 );
buf ( g4676 , g7 );
buf ( g4698 , g29 );
buf ( g4699 , g30 );
buf ( g4701 , g32 );
buf ( g4702 , g33 );
buf ( g4703 , g34 );
buf ( g4704 , g35 );
buf ( g4705 , g36 );
buf ( g4706 , g37 );
buf ( g4707 , g38 );
buf ( g4708 , g39 );
buf ( g4710 , g41 );
buf ( g4712 , g43 );
buf ( g4713 , g44 );
buf ( g4714 , g45 );
buf ( g4715 , g46 );
buf ( g4716 , g47 );
buf ( g4717 , g48 );
buf ( g4718 , g49 );
buf ( g4720 , g51 );
buf ( g4722 , g53 );
buf ( g4723 , g54 );
buf ( g4724 , g55 );
buf ( g4725 , g56 );
buf ( g4726 , g57 );
buf ( g4727 , g58 );
buf ( g4728 , g59 );
buf ( g4729 , g60 );
buf ( g4731 , g62 );
buf ( g4733 , g64 );
buf ( g4734 , g65 );
buf ( g4735 , g66 );
buf ( g4736 , g67 );
buf ( g4737 , g68 );
buf ( g4738 , g69 );
buf ( g4739 , g70 );
buf ( g4740 , g71 );
buf ( g4743 , g74 );
buf ( g4747 , g78 );
buf ( g4748 , g79 );
buf ( g4750 , g81 );
buf ( g4751 , g82 );
buf ( g4753 , g84 );
buf ( g4757 , g88 );
buf ( g4758 , g89 );
buf ( g4760 , g91 );
buf ( g4761 , g92 );
buf ( g4763 , g94 );
buf ( g4767 , g98 );
buf ( g4768 , g99 );
buf ( g4770 , g101 );
buf ( g4771 , g102 );
buf ( g4773 , g104 );
buf ( g4777 , g108 );
buf ( g4778 , g109 );
buf ( g4780 , g111 );
buf ( g4781 , g112 );
buf ( g4785 , g116 );
buf ( g4788 , g119 );
buf ( g4793 , g124 );
buf ( g4794 , g125 );
buf ( g4795 , g126 );
buf ( g4796 , g127 );
buf ( g4797 , g128 );
buf ( g4798 , g129 );
buf ( g4799 , g130 );
buf ( g4800 , g131 );
buf ( g4801 , g132 );
buf ( g4802 , g133 );
buf ( g4803 , g134 );
buf ( g4804 , g135 );
buf ( g4806 , g137 );
buf ( g4807 , g138 );
buf ( g4808 , g139 );
buf ( g4809 , g140 );
buf ( g4810 , g141 );
buf ( g4813 , g144 );
buf ( g4814 , g145 );
buf ( g4886 , g1377 );
nand ( g807 , g800 , g803 , g806 );
nand ( g653 , g645 , g647 , g650 , g652 );
nand ( g589 , g579 , g583 , g586 , g588 );
buf ( g975 , g543 );
not ( g1199 , g653 );
not ( g1245 , g807 );
nand ( g732 , g727 , g729 , g730 , g731 );
not ( g1135 , g525 );
nand ( g457 , g449 , g451 , g454 , g456 );
nand ( g1377 , g1363 , g1376 );
nand ( g446 , g4788 , g4785 );
not ( g447 , g4722 );
nor ( g448 , g446 , g447 );
not ( g449 , g448 );
not ( g450 , g4788 );
nand ( g451 , g450 , g4785 , g4701 );
not ( g452 , g4712 );
nor ( g453 , g452 , g4785 );
nand ( g454 , g453 , g4788 );
nor ( g455 , g4788 , g4785 );
nand ( g456 , g455 , g4733 );
not ( g466 , g4814 );
not ( g488 , g4814 );
nor ( g489 , g488 , g4813 );
not ( g495 , g4813 );
nor ( g501 , g4813 , g4814 );
not ( g511 , g4734 );
nor ( g512 , g511 , g4785 , g4788 );
nand ( g513 , g4788 , g4785 );
not ( g514 , g4723 );
nor ( g515 , g513 , g514 );
nor ( g516 , g512 , g515 );
not ( g517 , g516 );
not ( g518 , g4788 );
nand ( g519 , g518 , g4702 );
and ( g520 , g4785 , g519 );
not ( g521 , g4785 );
nand ( g522 , g4713 , g4788 );
and ( g523 , g521 , g522 );
nor ( g524 , g520 , g523 );
nor ( g525 , g517 , g524 );
not ( g534 , g4739 );
nor ( g535 , g534 , g4785 );
not ( g536 , g4788 );
nand ( g537 , g535 , g536 );
not ( g538 , g4788 );
nand ( g539 , g4785 , g538 , g4707 );
not ( g540 , g4785 );
nand ( g541 , g540 , g4788 , g4717 );
nand ( g542 , g4788 , g4728 , g4785 );
nand ( g543 , g537 , g539 , g541 , g542 );
not ( g550 , g4796 );
not ( g554 , g4813 );
not ( g555 , g4763 );
nand ( g556 , g554 , g555 , g4814 );
not ( g557 , g4753 );
nand ( g558 , g557 , g4813 , g4814 );
nor ( g559 , g4814 , g4743 );
nand ( g560 , g559 , g4813 );
not ( g561 , g4814 );
not ( g562 , g4773 );
nand ( g563 , g561 , g495 , g562 );
not ( g576 , g4785 );
nor ( g577 , g576 , g4788 );
not ( g578 , g4706 );
nand ( g579 , g577 , g578 );
not ( g580 , g4788 );
nor ( g581 , g580 , g4785 );
not ( g582 , g4716 );
nand ( g583 , g581 , g582 );
not ( g584 , g4738 );
nor ( g585 , g4785 , g4788 );
nand ( g586 , g584 , g585 );
not ( g587 , g4727 );
nand ( g588 , g587 , g4788 , g4785 );
nor ( g607 , g4814 , g4813 );
nand ( g608 , g607 , g4777 );
not ( g609 , g4814 );
nand ( g610 , g609 , g4747 , g4813 );
nand ( g611 , g608 , g610 );
not ( g625 , g4785 );
not ( g626 , g4731 );
not ( g627 , g4788 );
nand ( g628 , g625 , g626 , g627 );
not ( g629 , g4699 );
not ( g630 , g4788 );
nand ( g631 , g629 , g630 , g4785 );
not ( g632 , g4785 );
not ( g633 , g4710 );
nand ( g634 , g632 , g633 , g4788 );
not ( g635 , g4720 );
nand ( g636 , g635 , g4788 , g4785 );
nand ( g637 , g628 , g631 , g634 , g636 );
not ( g644 , g4715 );
nand ( g645 , g581 , g644 );
not ( g646 , g4705 );
nand ( g647 , g577 , g646 );
not ( g648 , g4737 );
nor ( g649 , g4785 , g4788 );
nand ( g650 , g648 , g649 );
not ( g651 , g4726 );
nand ( g652 , g651 , g4785 , g4788 );
not ( g658 , g4798 );
nor ( g666 , g4788 , g4740 );
not ( g667 , g4785 );
nand ( g668 , g666 , g667 );
not ( g669 , g4708 );
not ( g670 , g4788 );
nand ( g671 , g669 , g670 , g4785 );
not ( g672 , g4729 );
nand ( g673 , g672 , g4788 , g4785 );
not ( g674 , g4718 );
nand ( g675 , g667 , g674 , g4788 );
nand ( g676 , g668 , g671 , g673 , g675 );
not ( g677 , g676 );
not ( g678 , g677 );
not ( g685 , g4804 );
not ( g688 , g4761 );
nand ( g689 , g688 , g4813 , g4814 );
not ( g690 , g4771 );
nand ( g691 , g690 , g489 );
not ( g692 , g4781 );
nand ( g693 , g692 , g501 );
not ( g694 , g4751 );
nand ( g695 , g694 , g466 , g4813 );
not ( g704 , g4770 );
not ( g705 , g4814 );
nor ( g706 , g705 , g4813 );
nand ( g707 , g704 , g706 );
nor ( g708 , g4814 , g4750 );
nand ( g709 , g708 , g4813 );
not ( g710 , g4760 );
nand ( g711 , g710 , g4813 , g4814 );
not ( g712 , g4780 );
nor ( g713 , g4814 , g4813 );
nand ( g714 , g712 , g713 );
nand ( g715 , g707 , g709 , g711 , g714 );
not ( g720 , g4806 );
nand ( g725 , g4703 , g4785 );
nor ( g726 , g725 , g4788 );
not ( g727 , g726 );
not ( g728 , g4785 );
nand ( g729 , g728 , g4735 );
nand ( g730 , g728 , g4788 );
nand ( g731 , g4788 , g4724 );
not ( g739 , g4800 );
not ( g750 , g4807 );
not ( g771 , g4794 );
not ( g790 , g4810 );
nand ( g794 , g4788 , g4785 );
not ( g795 , g794 );
not ( g796 , g4725 );
and ( g797 , g795 , g796 );
nor ( g798 , g4788 , g4736 );
and ( g799 , g798 , g728 );
nor ( g800 , g797 , g799 );
not ( g801 , g4714 );
not ( g802 , g4785 );
nand ( g803 , g801 , g802 , g4788 );
not ( g804 , g4788 );
not ( g805 , g4704 );
nand ( g806 , g804 , g805 , g4785 );
not ( g813 , g4799 );
not ( g822 , g611 );
not ( g823 , g4813 );
nand ( g824 , g823 , g4767 , g4814 );
nand ( g825 , g4813 , g4757 , g4814 );
nand ( g826 , g824 , g825 , g4698 );
not ( g827 , g826 );
not ( g828 , g4748 );
nand ( g829 , g828 , g4813 );
not ( g830 , g4813 );
not ( g831 , g4778 );
nand ( g832 , g830 , g831 );
nor ( g833 , g4795 , g4814 );
nand ( g834 , g829 , g832 , g833 );
nor ( g835 , g4813 , g4768 );
not ( g836 , g835 );
not ( g837 , g4758 );
nand ( g838 , g837 , g4813 );
not ( g839 , g4795 );
nand ( g840 , g836 , g838 , g839 , g4814 );
nand ( g841 , g822 , g827 , g834 , g840 );
not ( g842 , g841 );
not ( g843 , g842 );
not ( g844 , g715 );
nand ( g845 , g844 , g4806 );
nand ( g846 , g4802 , g457 );
nand ( g847 , g560 , g563 );
not ( g848 , g847 );
not ( g849 , g556 );
not ( g850 , g849 );
nand ( g851 , g848 , g850 , g558 , g4803 );
nand ( g852 , g845 , g846 , g851 );
not ( g853 , g852 );
or ( g854 , g843 , g853 );
not ( g855 , g841 );
nand ( g856 , g689 , g693 );
not ( g857 , g856 );
and ( g858 , g691 , g695 );
nand ( g859 , g857 , g858 );
nor ( g860 , g859 , g685 );
nand ( g861 , g855 , g860 );
nand ( g862 , g854 , g861 );
not ( g863 , g862 );
buf ( g869 , g637 );
not ( g870 , g869 );
not ( g960 , g750 );
not ( g961 , g543 );
not ( g962 , g961 );
or ( g963 , g960 , g962 );
nand ( g964 , g963 , g4806 );
nor ( g965 , g611 , g826 );
nand ( g966 , g834 , g840 );
nand ( g967 , g965 , g966 );
not ( g968 , g967 );
or ( g969 , g961 , g678 );
nand ( g970 , g964 , g968 , g969 );
not ( g977 , g550 );
not ( g978 , g961 );
or ( g979 , g977 , g978 );
nand ( g980 , g979 , g4794 );
not ( g1005 , g4676 );
nand ( g1006 , g670 , g669 , g4785 );
not ( g1007 , g4729 );
nand ( g1008 , g1007 , g4788 , g4785 );
not ( g1009 , g4785 );
nand ( g1010 , g1009 , g674 , g4788 );
nand ( g1011 , g668 , g1006 , g1008 , g1010 );
nand ( g1134 , g4800 , g732 );
nand ( g1136 , g1135 , g4801 );
and ( g1137 , g1134 , g1136 );
nor ( g1138 , g1137 , g1005 );
not ( g1246 , g1245 );
not ( g1247 , g4809 );
nand ( g1248 , g965 , g966 );
not ( g1249 , g1248 );
not ( g1250 , g1249 );
or ( g1251 , g1247 , g1250 );
or ( g1252 , g658 , g1249 );
nand ( g1253 , g1251 , g1252 );
nand ( g1254 , g1253 , g1199 );
nor ( g1255 , g678 , g771 );
and ( g1256 , g859 , g685 );
buf ( g1257 , g715 );
and ( g1258 , g1257 , g720 );
nor ( g1259 , g1256 , g1258 );
not ( g1265 , g968 );
nand ( g1266 , g1265 , g980 , g969 );
nand ( g1267 , g1266 , g970 );
buf ( g1268 , g1248 );
or ( g1269 , g4801 , g1135 );
not ( g1270 , g732 );
nand ( g1271 , g1270 , g1136 , g739 );
nand ( g1272 , g1269 , g1271 );
nand ( g1273 , g1268 , g1138 );
nand ( g1274 , g813 , g1248 );
not ( g1275 , g1249 );
not ( g1276 , g790 );
or ( g1277 , g1275 , g1276 );
nand ( g1278 , g1277 , g1274 );
or ( g1279 , g1278 , g1246 );
nand ( g1280 , g1279 , g1254 );
nand ( g1281 , g863 , g1273 );
not ( g1282 , g4807 );
not ( g1283 , g968 );
or ( g1284 , g1282 , g1283 );
nand ( g1285 , g967 , g4796 );
nand ( g1286 , g1284 , g1285 );
not ( g1287 , g1011 );
nand ( g1288 , g1286 , g1287 );
and ( g1289 , g1267 , g1288 );
nor ( g1290 , g1249 , g1255 , g4793 );
not ( g1291 , g1290 );
not ( g1292 , g870 );
not ( g1293 , g1292 );
or ( g1294 , g1291 , g1293 );
and ( g1295 , g1287 , g4806 );
nor ( g1296 , g1295 , g4804 );
nand ( g1297 , g1292 , g1296 , g1249 );
nand ( g1298 , g1294 , g1297 );
nor ( g1299 , g1289 , g1298 );
not ( g1300 , g1286 );
buf ( g1301 , g975 );
not ( g1302 , g1301 );
or ( g1303 , g1300 , g1302 );
not ( g1304 , g4797 );
not ( g1305 , g1304 );
not ( g1306 , g1268 );
or ( g1307 , g1305 , g1306 );
not ( g1308 , g4808 );
nand ( g1309 , g1308 , g1249 );
nand ( g1310 , g1307 , g1309 );
buf ( g1311 , g589 );
or ( g1312 , g1310 , g1311 );
nand ( g1313 , g1303 , g1312 );
or ( g1314 , g1299 , g1313 );
not ( g1315 , g1253 );
nand ( g1316 , g4676 , g653 );
not ( g1317 , g1316 );
and ( g1318 , g1315 , g1317 );
and ( g1319 , g1310 , g1311 );
nor ( g1320 , g1318 , g1319 );
nand ( g1321 , g1314 , g1320 );
not ( g1326 , g457 );
nor ( g1327 , g4803 , g4802 );
nand ( g1328 , g1326 , g1327 );
not ( g1329 , g558 );
nor ( g1330 , g1329 , g847 , g849 );
and ( g1331 , g1328 , g1330 );
not ( g1332 , g4802 );
nand ( g1333 , g1332 , g1326 );
and ( g1334 , g1333 , g4803 );
nor ( g1335 , g1331 , g1334 );
nand ( g1349 , g1278 , g1273 , g807 );
and ( g1359 , g1280 , g4676 );
nor ( g1360 , g1359 , g1281 );
not ( g1361 , g1360 );
not ( g1362 , g1321 );
or ( g1363 , g1361 , g1362 );
not ( g1364 , g1268 );
not ( g1365 , g1272 );
or ( g1366 , g1364 , g1365 );
nand ( g1367 , g1366 , g1349 );
nor ( g1368 , g862 , g1005 );
and ( g1369 , g1367 , g1368 );
not ( g1370 , g861 );
not ( g1371 , g1335 );
or ( g1372 , g1370 , g1371 );
nand ( g1373 , g1372 , g1259 );
and ( g1374 , g842 , g845 );
and ( g1375 , g1373 , g1374 );
nor ( g1376 , g1369 , g1375 );
endmodule
